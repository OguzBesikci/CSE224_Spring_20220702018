magic
tech sky130A
magscale 1 2
timestamp 1745578439
<< nwell >>
rect 1066 2159 38862 37574
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 842 2128 38824 37584
<< obsm2 >>
rect 846 2139 38438 37573
<< metal3 >>
rect 0 37000 800 37120
rect 39200 37000 40000 37120
rect 0 32104 800 32224
rect 39200 32104 40000 32224
rect 0 27208 800 27328
rect 39200 27208 40000 27328
rect 0 22312 800 22432
rect 39200 22312 40000 22432
rect 0 17416 800 17536
rect 39200 17416 40000 17536
rect 0 12520 800 12640
rect 39200 12520 40000 12640
rect 0 7624 800 7744
rect 39200 7624 40000 7744
rect 0 2728 800 2848
rect 39200 2728 40000 2848
<< obsm3 >>
rect 798 37200 39200 37569
rect 880 36920 39120 37200
rect 798 32304 39200 36920
rect 880 32024 39120 32304
rect 798 27408 39200 32024
rect 880 27128 39120 27408
rect 798 22512 39200 27128
rect 880 22232 39120 22512
rect 798 17616 39200 22232
rect 880 17336 39120 17616
rect 798 12720 39200 17336
rect 880 12440 39120 12720
rect 798 7824 39200 12440
rect 880 7544 39120 7824
rect 798 2928 39200 7544
rect 880 2648 39120 2928
rect 798 2143 39200 2648
<< metal4 >>
rect 4208 2128 4528 37584
rect 4868 2128 5188 37584
rect 34928 2128 35248 37584
rect 35588 2128 35908 37584
<< metal5 >>
rect 1056 36642 38872 36962
rect 1056 35982 38872 36302
rect 1056 6006 38872 6326
rect 1056 5346 38872 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 38872 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 38872 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 38872 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 38872 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 37000 800 37120 6 in[0]
port 3 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 in[1]
port 4 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 in[2]
port 5 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 in[3]
port 6 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 in[4]
port 7 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 in[5]
port 8 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 in[6]
port 9 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 in[7]
port 10 nsew signal input
rlabel metal3 s 39200 37000 40000 37120 6 out[0]
port 11 nsew signal output
rlabel metal3 s 39200 32104 40000 32224 6 out[1]
port 12 nsew signal output
rlabel metal3 s 39200 27208 40000 27328 6 out[2]
port 13 nsew signal output
rlabel metal3 s 39200 22312 40000 22432 6 out[3]
port 14 nsew signal output
rlabel metal3 s 39200 17416 40000 17536 6 out[4]
port 15 nsew signal output
rlabel metal3 s 39200 12520 40000 12640 6 out[5]
port 16 nsew signal output
rlabel metal3 s 39200 7624 40000 7744 6 out[6]
port 17 nsew signal output
rlabel metal3 s 39200 2728 40000 2848 6 out[7]
port 18 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 567068
string GDS_FILE /openlane/designs/twos_complement/runs/RUN_2025.04.25_10.53.07/results/signoff/twos_complement.magic.gds
string GDS_START 92926
<< end >>

